`timescale 1ns/1ps // Compiler directive: sets the time unit to 1ns and precision to 1ps for simulation.

module eSPI_Master #( // Defines the start of a module named 'eSPI_Master'. '#' begins the parameter list.
    parameter DATA_WIDTH = 8, // Defines a configurable parameter 'DATA_WIDTH' with a default value of 8.
    parameter CLK_DIVISOR = 4 // Defines a parameter 'CLK_DIVISOR' for the sclk generator, default is 4.
  ) ( // Begins the list of module ports (inputs and outputs).
    input  logic clk, // Input port: 'clk', the main system clock. 'logic' is a 4-state data type.
    input  logic reset_n, // Input port: 'reset_n', an active-low asynchronous reset. The '_n' denotes active-low.

    // Host interface // Comment: The following ports connect to the host system.
    input  logic start_transaction, // Input port: A signal from the host to initiate a transaction.
    input  logic [7:0] command, // Input port: An 8-bit command value from the host.
    input  logic [DATA_WIDTH-1:0] write_data, // Input port: Data to be written, width is parameterized by DATA_WIDTH.
    output logic [DATA_WIDTH-1:0] read_data, // Output port: Data read from the slave, width is parameterized.
    output logic transaction_done, // Output port: A flag indicating the transaction has finished.

    // eSPI physical signals // Comment: The following ports connect to the physical eSPI bus.
    output logic sclk, // Output port: The eSPI serial clock, generated by this master module.
    output logic cs_n, // Output port: The active-low chip select signal for the eSPI slave.
    inout  wire io0 // Bidirectional port: The main data line (io0). 'inout' for bidirectional, 'wire' for physical connection.
  ); // Ends the port list.

  // FSM state definitions // Comment: Defines the states for the Finite State Machine (FSM).
  typedef enum logic [1:0] { // 'typedef enum' creates a custom data type for the FSM states, using 2 bits.
            IDLE, // State: Waiting for a transaction to start.
            COMMAND_PHASE, // State: Sending the 8-bit command to the slave.
            TAR_PHASE, // State: Turn-Around-Time phase, bus direction changes from master-drive to slave-drive.
            RESPONSE_PHASE // State: Master receives data from the slave.
          } state_t; // Names the new enumerated type 'state_t'.

  state_t current_state, next_state; // Declares two signals of type 'state_t' to hold the FSM's current and next state.

  // Internal registers and signals // Comment: Declaration of internal signals and registers used within the module.
  logic [7:0] command_reg; // An 8-bit register to store the command for the transaction's duration.
  logic [DATA_WIDTH-1:0] read_data_reg; // A register to capture incoming data from the slave.
  logic [DATA_WIDTH-1:0] write_data_reg; // A register to store the outgoing data to be written.
  logic [$clog2(DATA_WIDTH)-1:0] bit_counter; // A counter for tracking bits. Width is calculated by '$clog2' to be just large enough for DATA_WIDTH.
  logic clk_enable; // A control signal to enable the 'sclk' generator only during a transaction.
  logic [$clog2(CLK_DIVISOR)-1:0] clk_div_counter; // A counter for the clock divider. Width is calculated by '$clog2'.
  logic sclk_d; // A delayed version of 'sclk' (d for delay), used for edge detection.
  logic sclk_negedge; // A pulse signal that goes high for one 'clk' cycle on the falling edge of 'sclk'.

  // Tri-state driver for io0 // Comment: Logic for the bidirectional 'io0' pin.
  logic io0_o; // The output value to drive onto 'io0' when the master is transmitting.
  logic io0_t; // The tri-state enable signal. '1' = high-impedance (input), '0' = drive 'io0_o' (output).
  assign io0 = (io0_t) ? 1'bz : io0_o; // 'assign' creates a continuous assignment. If 'io0_t' is true, 'io0' is high-impedance ('1'bz'); otherwise, it's driven by 'io0_o'.

  // Clock divider for SCLK generation // Comment: This block generates the eSPI clock ('sclk') from the system clock ('clk').
  always_ff @(posedge clk or negedge reset_n) // 'always_ff' describes sequential logic (flip-flops). It triggers on the 'posedge' (rising edge) of 'clk' or 'negedge' (falling edge) of 'reset_n'.
  begin // Starts the procedural block.
    if (!reset_n) // Checks for the active-low asynchronous reset condition. '!' is the logical NOT operator.
    begin // Starts the reset logic block.
      clk_div_counter <= 0; // On reset, asynchronously set the clock divider counter to 0. '<=' is the non-blocking assignment for sequential logic.
      sclk <= 0; // On reset, asynchronously set the 'sclk' output to 0.
    end // Ends the reset logic block.
    else if (clk_enable) // If not in reset, this logic is evaluated on 'posedge clk'. Checks if clock generation is enabled.
    begin // Starts the enabled clock divider logic.
      if (clk_div_counter == CLK_DIVISOR-1) // Checks if the counter has reached its maximum value.
      begin // Starts the counter wrap-around logic.
        clk_div_counter <= 0; // Resets the counter back to 0.
        sclk <= ~sclk; // Toggles the 'sclk' signal. '~' is the bitwise NOT operator, flipping the bit.
      end // Ends the counter wrap-around logic.
      else // If the counter has not reached its max value.
      begin // Starts the counter increment logic.
        clk_div_counter <= clk_div_counter + 1; // Increments the counter by 1.
      end // Ends the counter increment logic.
    end // Ends the enabled clock divider logic.
    else // If clock generation is not enabled (e.g., in IDLE state).
    begin // Starts the disabled clock divider logic.
      clk_div_counter <= 0; // Keeps the counter at 0.
      sclk <= 0; // Keeps the 'sclk' output low.
    end // Ends the disabled clock divider logic.
  end // Ends the 'always_ff' block.

  // SCLK edge detection in clk domain // Comment: This logic detects the falling edge of 'sclk' and creates a single-cycle pulse.
  always_ff @(posedge clk or negedge reset_n) // A sequential block, sensitive to the system clock and reset.
  begin // Starts the block.
    if (!reset_n) // Asynchronous reset condition.
    begin // Starts reset logic.
      sclk_d <= 1'b0; // On reset, set the delayed sclk signal to 0. '1'b0' is a 1-bit binary value of 0.
    end // Ends reset logic.
    else // Synchronous part, on the 'posedge clk'.
    begin // Starts synchronous logic.
      sclk_d <= sclk; // On each clock edge, sample the current value of 'sclk' into 'sclk_d', creating a one-cycle delay.
    end // Ends synchronous logic.
  end // Ends the 'always_ff' block.
  assign sclk_negedge = sclk_d & ~sclk; // Continuous assignment. 'sclk_negedge' is high only when the previous value ('sclk_d') was 1 and the current value ('sclk') is 0. '&' is the bitwise AND.

  // FSM sequential block // Comment: This is the main sequential block for the FSM state and other registers.
  always_ff @(posedge clk or negedge reset_n) // This block describes all the registers that change on the clock edge.
  begin // Starts the block.
    if (!reset_n) // Asynchronous reset condition.
    begin // Starts reset logic.
      current_state    <= IDLE; // Resets the FSM to the IDLE state.
      bit_counter      <= 0; // Resets the bit counter.
      cs_n             <= 1; // De-asserts the chip select signal (active low, so 1 is inactive).
      io0_t            <= 1; // Puts the 'io0' line in high-impedance (tri-state) mode.
      read_data_reg    <= 0; // Clears the read data register.
      transaction_done <= 0; // Clears the transaction done flag.
    end // Ends reset logic.
    else // Synchronous part, on the 'posedge clk'.
    begin // Starts synchronous logic.
      current_state    <= next_state; // Updates the current state with the value calculated in the combinational 'always_comb' block.
      transaction_done <= 0; // Default assignment: clears 'transaction_done' on every clock cycle unless set otherwise.

      case (current_state) // 'case' statement to describe behavior based on the 'current_state'.
        IDLE: // Behavior for the IDLE state.
        begin // Starts IDLE state logic.
          if (start_transaction) // Checks if a new transaction is requested by the host.
          begin // Starts transaction initiation logic.
            command_reg    <= command; // Latches the command from the host interface into an internal register.
            write_data_reg <= write_data; // Latches the write data from the host interface.
            cs_n           <= 0; // Asserts the chip select signal (drives it low).
            io0_t          <= 0; // Enables the output driver for 'io0' (stops tri-stating).
            bit_counter    <= 0; // Resets the bit counter for the new transaction.
          end // Ends transaction initiation logic.
        end // Ends IDLE state logic.

        COMMAND_PHASE: // Behavior for the COMMAND_PHASE state.
        begin // Starts COMMAND_PHASE logic.
          // Slave samples on posedge sclk, so we change our output on the negedge of sclk for better timing margin.
          if (sclk_negedge) // Checks for the single-cycle pulse indicating a falling edge on 'sclk'.
          begin // Starts bit transmission logic.
            io0_o <= command_reg[7-bit_counter]; // Drives the next bit of the command onto the 'io0' line.
            if (bit_counter == 7) // Checks if all 8 bits of the command have been sent.
            begin // Starts logic for the last bit.
              io0_t <= 1; // Tri-state the bus in preparation for the Turn-Around phase.
            end // Ends logic for the last bit.
            else // If not the last bit.
            begin // Starts bit counter increment logic.
              bit_counter <= bit_counter + 1; // Increments the bit counter to send the next bit.
            end // Ends bit counter increment logic.
          end // Ends bit transmission logic.
        end // Ends COMMAND_PHASE logic.

        TAR_PHASE: // Behavior for the Turn-Around-Time phase.
        begin // Starts TAR_PHASE logic.
          // This phase is for bus direction change. We reset the bit counter for the next phase.
          bit_counter <= 0; // Resets the bit counter to prepare for the RESPONSE_PHASE.
        end // Ends TAR_PHASE logic.

        RESPONSE_PHASE: // Behavior for the RESPONSE_PHASE state.
        begin // Starts RESPONSE_PHASE logic.
          // Slave drives on posedge sclk, so we sample on negedge sclk for better timing margin.
          if (sclk_negedge) // Checks for the falling edge of 'sclk' to sample the incoming data.
          begin // Starts bit reception logic.
            read_data_reg[DATA_WIDTH-1-bit_counter] <= io0; // Samples the 'io0' line and stores the bit in the read data register.
            if (bit_counter == DATA_WIDTH-1) // Checks if all bits of the response have been received.
            begin // Starts logic for the last bit.
              cs_n             <= 1; // De-asserts chip select to end the transaction.
              transaction_done <= 1; // Sets the flag to signal the host that the transaction is complete.
            end // Ends logic for the last bit.
            else // If not the last bit.
            begin // Starts bit counter increment logic.
              bit_counter <= bit_counter + 1; // Increments the bit counter to receive the next bit.
            end // Ends bit counter increment logic.
          end // Ends bit reception logic.
        end // Ends RESPONSE_PHASE logic.
      endcase // Ends the 'case' statement for the FSM states.
    end // Ends the synchronous logic block.
  end // Ends the 'always_ff' block.

  // Next-state logic and outputs // Comment: This block describes the combinational logic for FSM state transitions and outputs.
  always_comb // 'always_comb' declares that the logic inside is purely combinational. The block re-evaluates whenever any input signal changes.
  begin // Starts the combinational block.
    next_state = current_state; // Default assignment: the next state is the same as the current state unless a transition condition is met.
    clk_enable = (current_state != IDLE); // The 'sclk' generator is enabled in any state except IDLE.
    read_data  = read_data_reg; // The module's output 'read_data' is continuously driven by the internal 'read_data_reg'.

    case (current_state) // 'case' statement to determine the next state based on the current state and inputs.
      IDLE: // Transition logic for the IDLE state.
      begin // Starts IDLE transition logic.
        if (start_transaction) // If a transaction is requested.
          next_state = COMMAND_PHASE; // Transition to the COMMAND_PHASE.
      end // Ends IDLE transition logic.

      COMMAND_PHASE: // Transition logic for the COMMAND_PHASE state.
      begin // Starts COMMAND_PHASE transition logic.
        if (sclk_negedge && bit_counter == 7) // If the last bit of the command has just been sent.
          next_state = TAR_PHASE; // Transition to the TAR_PHASE.
      end // Ends COMMAND_PHASE transition logic.

      TAR_PHASE: // Transition logic for the TAR_PHASE state.
      begin // Starts TAR_PHASE transition logic.
        // This is a single-cycle state to allow for bus turn-around.
        next_state = RESPONSE_PHASE; // Unconditionally transition to the RESPONSE_PHASE on the next clock cycle.
      end // Ends TAR_PHASE transition logic.

      RESPONSE_PHASE: // Transition logic for the RESPONSE_PHASE state.
      begin // Starts RESPONSE_PHASE transition logic.
        if (sclk_negedge && bit_counter == DATA_WIDTH-1) // If the last bit of the response has just been received.
          next_state = IDLE; // Transition back to the IDLE state.
      end // Ends RESPONSE_PHASE transition logic.
    endcase // Ends the 'case' statement for state transitions.
  end // Ends the 'always_comb' block.

endmodule // Ends the module definition.

